`timescale 1ns / 1ps
 
module InstructionDecode(Clk, Rst, Instruction, WriteData, WriteRegister);

   // Inputs   
   input Clk, Rst;
   input [31:0] Instruction;
   input [31:0] WriteData;
   input [4:0] WriteRegister;
   
   // Outputs
   output ReadData1, ReadData2;
   
   // Control Signals
   
   
   
   
   
endmodule