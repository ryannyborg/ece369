`timescale 1ns / 1ps
 
module WriteBack(Clk, Rst);
   
   input Clk, Rst;
   
   
   
   
endmodule