`timescale 1ns / 1ps

module ShiftLeft2_tb();

    ShiftLeft2 u0(
    
    );
    

endmodule
