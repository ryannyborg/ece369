`timescale 1ns / 1ps
 
module Memory(Clk, Rst);
   
   input Clk, Rst;
   
   
   
   
endmodule