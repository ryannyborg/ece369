`timescale 1ns / 1ps
 
module TopLevel(Clk, Rst);
   
   input Clk, Rst;
   
   
   
   
endmodule