`timescale 1ns / 1ps
 
module Execution(Clk, Rst);
   
   input Clk, Rst;
   
   
   
   
endmodule