`timescale 1ns / 1ps

module EXAdder_tb();

    EXAdder u0(
        
    );

endmodule
