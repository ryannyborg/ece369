`timescale 1ns / 1ps

module IFIDRegister_tb();
    
    IFIDRegister u0(
    
    );
    
endmodule
